library verilog;
use verilog.vl_types.all;
entity timer_1ms_vlg_vec_tst is
end timer_1ms_vlg_vec_tst;
