library verilog;
use verilog.vl_types.all;
entity Tempo_umMs_vlg_check_tst is
    port(
        clk_umMs        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Tempo_umMs_vlg_check_tst;
