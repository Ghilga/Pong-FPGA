library verilog;
use verilog.vl_types.all;
entity Tempo_umMs_vlg_vec_tst is
end Tempo_umMs_vlg_vec_tst;
