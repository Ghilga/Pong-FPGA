library verilog;
use verilog.vl_types.all;
entity clk_pixel_vlg_vec_tst is
end clk_pixel_vlg_vec_tst;
