library verilog;
use verilog.vl_types.all;
entity clk_pixel_vlg_check_tst is
    port(
        clk_pixel       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end clk_pixel_vlg_check_tst;
